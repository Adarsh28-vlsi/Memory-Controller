`timescale 1ns / 1ps
module controller #(
  parameter R = 4,
  parameter C = 4,
  parameter N = 4
)(
  input wire clk,
  input wire rst,
  input wire cs,
  input wire req,
  input wire rw,
  input wire [$clog2(R*C)-1:0] addr,
  input wire valid,
  output reg ready,
  output wire [$clog2(R)-1:0] ar,
  output wire [$clog2(C)-1:0] ac
);
  assign ar = addr[$clog2(R*C)-1 -: $clog2(R)];
  assign ac = addr[$clog2(C)-1:0];
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      ready <= 1'b0;
    end else begin
      if (cs) begin
        if (req && !rw)
          ready <= 1'b1;
        else if (valid)
          ready <= 1'b1;
        else
          ready <= 1'b0;
      end else begin
        ready <= 1'b0;
      end
    end
  end
endmodule
