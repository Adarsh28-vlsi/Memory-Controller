`timescale 1ns / 1ps
module tb_sp;
  parameter R = 4;
  parameter C = 4;
  parameter N = 4;
  reg clk = 0;
  reg rst = 1;
  reg cs = 0, req = 0, rw = 0;
  reg [$clog2(R*C)-1:0] addr = 0;
  reg [N-1:0] Qi = 0;
  wire [N-1:0] Qa;
  wire valid, ready;
  top_module #(.R(R), .C(C), .N(N)) dut (
    .clk(clk), .rst(rst), .cs(cs),
    .req(req), .rw(rw), .addr(addr),
    .Qi(Qi), .Qa(Qa), .valid(valid), .ready(ready)
  );
  always #5 clk = ~clk;
  initial #25 rst = 0;
  initial begin
    @(negedge rst);
    cs = 1; addr = 4'd3; Qi = 4'h01; rw = 0; req = 1;
    @(posedge clk);
    req = 1; @(posedge clk);
    cs = 1; addr = 4'd3; rw = 1; req = 1;
    @(posedge clk);
    cs = 1; addr = 4'd5; Qi = 4'd06; rw = 0; req = 1;
    @(posedge clk);

    @(posedge clk);
    req = 1; @(posedge clk);
    cs = 1; addr = 4'd5; rw = 1; req = 1;
    @(posedge clk);
    $finish;
  end
endmodule
